module xor_op (
	input a1,
	input a2,
	output c
);

	assign c = a1^a2;

endmodule