module and_op (
	a1,
	a2,
	c
);

input a1,a2;
output c;


	assign c = a1 & a2;

endmodule