module not_op (
	input a,
	output c
);

	assign c = ~a;

endmodule